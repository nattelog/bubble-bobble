nattelog@c-213-14.eduroam.liu.se.70510