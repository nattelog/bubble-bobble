-- The CPU

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity cpu is
    Port (clk,rst : in  STD_LOGIC);
end cpu;

architecture behavioral of cpu is
  signal buss : STD_LOGIC_VECTOR(2 downto 0);
begin

-- ** ASR **

-- ** Programminne **

-- ** IR **

-- ** K1 **

-- ** K2 **

-- ** µPC **

-- ** µM **

-- ** Flaggor (Z, N, C, O, L)

-- ** GR **

-- ** RP (registerpekare) **

-- ** ALU **

-- ** AR **

-- ** PC **

end behavioral;
