nattelog@c-213-129.eduroam.liu.se.5058