-- The CPU

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity cpu is
    Port ( clk,rst : in  STD_LOGIC
    );
end cpu;

architecture behavioral of cpu is
begin

end behavioral;