nattelog@natanaels-mbp.mynet.73264