nattelog@localhost.221