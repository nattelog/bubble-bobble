-- The CPU
-- This architecture follows the same architecture as in
-- Lab 1 in the course TSEA83, except for some modifications.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity cpu is
  Port (clk,rst : in  STD_LOGIC);
end cpu;

architecture behavioral of cpu is

  -- Main registers for the CPU
  signal BUSS, IR, PM, PC, AR, GRx : STD_LOGIC_VECTOR(31 downto 0);

  -- Control-unit
  signal controlword : STD_LOGIC_VECTOR(0 to 23);
  signal mPC : STD_LOGIC_VECTOR(6 downto 0);
  type mM is array(0 to 127) of controlword;
  type kM is array(0 to 15) of STD_LOGIC_VECTOR(6 downto 0); -- K-registers
  type gR is array(0 to 15) of STD_LOGIC_VECTOR(31 downto 0); -- General registers

  -- Memory-unit
  signal programword : STD_LOGIC_VECTOR(31 downto 0);
  type pM is array(0 to 65535) of programword;

  -- Signals from controlword
  alias alu : STD_LOGIC_VECTOR(3 downto 0) is controlword(0 to 3);
  alias tb : STD_LOGIC_VECTOR(2 downto 0) is controlword(4 to 6);
  alias fb : STD_LOGIC_VECTOR(2 downto 0) is controlword(7 to 9);
  alias p : STD_LOGIC is controlword(10);
  alias lc : STD_LOGIC_VECTOR(1 downto 0) is controlword(11 to 12);
  alias seq : STD_LOGIC_VECTOR(3 downto 0) is controlword(13 to 16);
  alias madr : STD_LOGIC_VECTOR(6 downto 0) is controlword(17 to 23);

  -- Signals from programword
  alias op : STD_LOGIC_VECTOR(3 downto 0) is programword(31 downto 28);
  alias grx : STD_LOGIC_VECTOR(3 downto 0) is programword(27 downto 24);
  alias m : STD_LOGIC_VECTOR(1 downto 0) is programword(23 downto 22);
  alias padr : STD_LOGIC_VECTOR(15 downto 0) is programword(15 downto 0);

  -- K1
  constant K1 : kM := (
    X"00",      -- 0x0 : LDA
    X"00",      -- 0x1 : STR
    X"00",      -- 0x2 : ADD
    X"00",      -- 0x3 : SUB
    X"00",      -- 0x4 : CMP
    X"00",      -- 0x5 : AND
    X"00",      -- 0x6 : OR
    X"00",      -- 0x7 : LSR
    X"00",      -- 0x8 : LSL
    X"00",      -- 0x9 : BRA
    X"00",      -- 0xa : BRG
    X"00",      -- 0xb : BNE
    X"00",      -- 0xc : BRE
    X"00",      -- 0xd : BRC
    X"00",      -- 0xe : JSR
    X"00"       -- 0xf : RTS
    );

  -- K2
  constant K2 : kM := (
    X"00",      -- 0x0 : Direct
    X"00",      -- 0x1 : Constant
    X"00",      -- 0x2 : Indirect
    X"00",      -- 0x3 : Indexed
    others => X"00"
    );

  -- Micromemory
  constant mMem : mM := (
    others => X"00"
    );

  -- Programmemory
  signal pMem : pM := (
    others => X"00"
    );     
  
begin

  -- ** BUSS  **

  process (clk)
  begin
    if rising_edge(clk) then
      if (rst = '1') then
        BUSS <= (others => '0');
      end if;
    end if;
  end process;

  -- to bus
  case tb is

    -- read from IR
    when "001" =>
      BUSS <= IR;

    -- read from PM
    when "010" =>
      BUSS <= PM;

    -- read from PC 
    when "011" =>
      BUSS <= PC;

    -- read from AR  
    when "100" =>
      BUSS <= AR;

    -- read from GRx
    when "110" =>
      BUSS <= GRx;

    -- do nothing
    when others =>
      
  end case;

  -- from bus
  case fb is

    -- write to IR
    when "001" =>
      IR <= BUSS;

    -- write to PM
    when "010" =>
      PM <= BUSS;

    -- write to PC
    when "011" =>
      PC <= BUSS;

    -- write to GRx
    when "110" =>
      GRx <= BUSS;

    -- write to ASR
    when "111" =>
      ASR <= BUSS;

    -- do nothing
    when others =>  
    
  end case;

  -- ** Micromemory **

  process (clk)
  begin
    if rising_edge(clk) then
      if (rst = '1') then
        mPC <= (others => '0');
        controlword <= (others => '0');

      else
        controlword <= mMem(CONV_INTEGER(mPC));
        
      end if;
    end if;
  end process;
  
  -- ** ASR **

  process (clk)
  begin
    if rising_edge(clk) then
      if (rst = '1') then
        ASR <= (others => '0');

      elsif (fb = "111")
        
        
      end if;
    end if;
  end process;

  -- ** Programmemory **

  -- ** IR **

  -- ** µPC **

  -- ** SuPC

  -- ** Flaggor (Z, N, C, O, L)

  -- ** GR **

  -- ** RP (registerpekare) **

  -- ** ALU **

  -- ** AR **

  -- ** PC **

end behavioral;
